module telegram

pub struct WebAppInfo {
	url string [required] // 	An HTTPS URL of a Web App to be opened with additional data as specified in Initializing Web Apps
}
