module telegram

pub struct ChatMemberUpdated {
}
