module telegram

struct GeneralForumTopicHidden {

}
