module main

import telegram

fn main() {
	println('Hello World!')
}
