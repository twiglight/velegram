module telegram

pub struct VideoChatStarted {
}
