module telegram

struct ChatMemberUpdated {

}
