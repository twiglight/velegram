module telegram

pub struct ForumTopicReopened {
}
