module telegram

pub struct ForumTopicClosed {
}
