module telegram
