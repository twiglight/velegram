module telegram

pub struct GeneralForumTopicUnhidden {
}
