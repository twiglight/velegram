module telegram

struct WriteAccessAllowed {

}
