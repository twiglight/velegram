module telegram

struct ForumTopicReopened {

}
