module telegram

pub struct ChatJoinRequest {
}
