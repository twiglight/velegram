module telegram

struct GeneralForumTopicUnhidden {

}
