module telegram

pub struct VideoChatScheduled {
	start_date int [required] // 	Point in time (Unix timestamp) when the video chat is supposed to be started by a chat administrator
}
