module telegram

pub struct WriteAccessAllowed {
}
