module telegram

pub struct GeneralForumTopicHidden {
}
