module telegram

struct ChatJoinRequest {

}
