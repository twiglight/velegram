module telegram

struct VideoChatStarted {

}
