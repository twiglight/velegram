module telegram

struct VideoChatEnded {
	duration int [required] 			// 	Video chat duration in seconds
}
