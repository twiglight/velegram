module telegram

struct ForumTopicClosed {
	
}
